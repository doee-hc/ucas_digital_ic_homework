// Component Name   : sqrt_u32
// Component Version: 
// Release Type     : 
//  ------------------------------------------------------------------------

// 
// Release version :  
// File Version    :  
// Revision: 
//
//
// File    : design/sqrt_u32/rtl/sqrt_u32.v
// Author  : Huhc
// Date    : 2023-12-28 20:41:45
// Abstract: 
module sqrt_u32(

);


endmodule

